//=======================================================
//  This is the top level file
//=======================================================

// This code is implements a BCD to 7-Segment Decoder using verilog
// We have used Hierarchical Design to implement our circuit
// This is the top level file
// The bcd7segment module is initialized by giving the proper signals
// All the deductions for the 7-segment display segments can be read on the link below
// https://www.focuslk.com/design-of-bcd-to-7-segment-display-decoder-using-logic-gates/



//=======================================================
//  This code is generated by Terasic System Builder
//=======================================================

module DE10_LITE_TOP(

	//////////// CLOCK //////////
	input 		          		ADC_CLK_10,
	input 		          		MAX10_CLK1_50,
	input 		          		MAX10_CLK2_50,

	//////////// SDRAM //////////
	output		    [12:0]		DRAM_ADDR,
	output		     [1:0]		DRAM_BA,
	output		          		DRAM_CAS_N,
	output		          		DRAM_CKE,
	output		          		DRAM_CLK,
	output		          		DRAM_CS_N,
	inout 		    [15:0]		DRAM_DQ,
	output		          		DRAM_LDQM,
	output		          		DRAM_RAS_N,
	output		          		DRAM_UDQM,
	output		          		DRAM_WE_N,

	//////////// SEG7 //////////
	output		     [7:0]		HEX0,
	output		     [7:0]		HEX1,
	output		     [7:0]		HEX2,
	output		     [7:0]		HEX3,
	output		     [7:0]		HEX4,
	output		     [7:0]		HEX5,

	//////////// KEY //////////
	input 		     [1:0]		KEY,

	//////////// LED //////////
	output		     [9:0]		LEDR,

	//////////// SW //////////
	input 		     [9:0]		SW,

	//////////// VGA //////////
	output		     [3:0]		VGA_B,
	output		     [3:0]		VGA_G,
	output		          		VGA_HS,
	output		     [3:0]		VGA_R,
	output		          		VGA_VS,

	//////////// Accelerometer //////////
	output		          		GSENSOR_CS_N,
	input 		     [2:1]		GSENSOR_INT,
	output		          		GSENSOR_SCLK,
	inout 		          		GSENSOR_SDI,
	inout 		          		GSENSOR_SDO,

	//////////// Arduino //////////
	inout 		    [15:0]		ARDUINO_IO,
	inout 		          		ARDUINO_RESET_N
);



//=======================================================
//  REG/WIRE declarations
//=======================================================




//=======================================================
//  Structural coding
//=======================================================

//we need 4 inputs as the BCD - We take switches 0 to 4 in our Terrasic DE-10 lite
//we need 8 bit output for the display - We select Hex display 0 as out diplay
	
bcd7segment bcdCircuit(SW[3:0],HEX0);  //Making an instance of the BCD to 7 segment decoder
	
//uncomment this to run the circuit using behavioral modelling
//bcd7segmentBehavioral bcdCircuit1(SW[3:0],HEX0); //Making an instance of the BCD to 7 segment decoder




endmodule
